package ahb2apb_test_pkg;

	import uvm_pkg::*;
//include uvm_macros.sv
`include "uvm_macros.svh"
`include "write_xtn.sv"
`include "ahb2apb_master_agent_config.sv"
`include "ahb2apb_slave_agent_config.sv"
`include "ahb2apb_env_config.sv"
`include "ahb2apb_master_driver.sv"
`include "ahb2apb_master_monitor.sv"
`include "ahb2apb_master_sequencer.sv"
`include "ahb2apb_master_agent.sv"
`include "ahb2apb_master_agt_top.sv"
`include "ahb2apb_master_sequence.sv"


`include "read_xtn.sv"
`include "ahb2apb_slave_monitor.sv"
`include "ahb2apb_slave_sequencer.sv"
`include "ahb2apb_slave_sequence.sv"
`include "ahb2apb_slave_driver.sv"
`include "ahb2apb_slave_agent.sv"
`include "ahb2apb_slave_agt_top.sv"

`include "ahb2apb_virtual_sequencer.sv"
`include "ahb2apb_virtual_sequences.sv"
`include "ahb2apb_scoreboard.sv"

`include "ahb2apb_env.sv"

`include "ahb2apb_testcases.sv"
endpackage
